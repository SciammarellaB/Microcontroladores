CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
290 50 30 200 9
38 98 1498 837
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 98 1498 837
143654930 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 810 178 0 1 11
0 6
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V14
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 779 215 0 1 11
0 7
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V13
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 676 99 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V12
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 650 99 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 625 99 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 599 99 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 391 369 0 1 11
0 12
0
0 0 21360 0
2 0V
-33 -4 -19 4
2 V8
-33 -14 -19 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 391 345 0 1 11
0 13
0
0 0 21360 0
2 0V
-33 -4 -19 4
2 V7
-33 -14 -19 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 391 322 0 1 11
0 14
0
0 0 21360 0
2 0V
-33 -4 -19 4
2 V6
-33 -14 -19 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 391 298 0 1 11
0 15
0
0 0 21360 0
2 0V
-33 -4 -19 4
2 V5
-33 -14 -19 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 392 213 0 1 11
0 17
0
0 0 21360 0
2 0V
-33 -2 -19 6
2 V3
-33 -14 -19 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 392 239 0 1 11
0 16
0
0 0 21360 0
2 0V
-34 -1 -20 7
2 V4
-34 -14 -20 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 392 187 0 1 11
0 18
0
0 0 21360 0
2 0V
-33 -2 -19 6
2 V2
-32 -14 -18 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3834 0 0
0
0
13 Logic Switch~
5 392 161 0 1 11
0 19
0
0 0 21360 0
2 0V
-33 -4 -19 4
2 V1
-33 -14 -19 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3363 0 0
0
0
4 LED~
171 959 257 0 1 2
10 5
0
0 0 368 0
1 P
-4 13 3 21
2 D8
-7 24 7 32
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
7668 0 0
0
0
4 LED~
171 925 257 0 1 2
10 4
0
0 0 368 0
1 G
-4 13 3 21
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4718 0 0
0
0
4 LED~
171 892 257 0 1 2
10 3
0
0 0 368 0
3 A=B
-11 13 10 21
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3874 0 0
0
0
4 LED~
171 861 257 0 1 2
10 2
0
0 0 368 0
4 Cn 4
-14 13 14 21
0
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
6671 0 0
0
0
4 LED~
171 798 311 0 1 2
10 23
0
0 0 880 0
4 LED1
-14 13 14 21
2 D4
-7 24 7 32
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3789 0 0
0
0
4 LED~
171 765 311 0 1 2
10 22
0
0 0 880 0
4 LED1
-14 13 14 21
2 D3
-7 24 7 32
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4871 0 0
0
0
4 LED~
171 733 311 0 1 2
10 21
0
0 0 880 0
4 LED1
-14 13 14 21
2 D2
-7 24 7 32
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3750 0 0
0
0
4 LED~
171 700 311 0 1 2
10 20
0
0 0 880 0
4 LED1
-14 13 14 21
2 D1
-7 24 7 32
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
8778 0 0
0
0
7 74LS181
132 640 233 0 22 45
0 8 9 10 11 19 18 17 16 15
14 13 12 6 7 2 3 4 5 20
21 22 23
0
0 0 13040 0
7 74LS181
-24 -69 25 -61
2 U1
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 0 1 0 0 0
1 U
538 0 0
0
0
22
15 1 2 0 0 4224 0 23 18 0 0 5
672 224
816 224
816 217
861 217
861 247
16 1 3 0 0 4224 0 23 17 0 0 5
672 233
823 233
823 225
892 225
892 247
17 1 4 0 0 4224 0 23 16 0 0 5
678 242
832 242
832 232
925 232
925 247
18 1 5 0 0 4224 0 23 15 0 0 5
678 251
840 251
840 239
959 239
959 247
13 1 6 0 0 4224 0 23 1 0 0 4
672 188
741 188
741 178
796 178
14 1 7 0 0 4224 0 23 2 0 0 4
672 197
727 197
727 215
765 215
1 1 8 0 0 8320 0 23 6 0 0 5
608 188
573 188
573 131
599 131
599 111
2 1 9 0 0 8320 0 23 5 0 0 5
608 197
579 197
579 141
625 141
625 111
3 1 10 0 0 12416 0 23 4 0 0 5
608 206
588 206
588 151
650 151
650 111
4 1 11 0 0 12416 0 23 3 0 0 5
608 215
597 215
597 160
676 160
676 111
1 12 12 0 0 12416 0 7 23 0 0 4
403 369
502 369
502 287
602 287
1 11 13 0 0 4224 0 8 23 0 0 4
403 345
518 345
518 278
602 278
1 10 14 0 0 4224 0 9 23 0 0 4
403 322
537 322
537 269
602 269
1 9 15 0 0 4224 0 10 23 0 0 4
403 298
556 298
556 260
602 260
1 8 16 0 0 12416 0 12 23 0 0 4
404 239
502 239
502 251
602 251
1 7 17 0 0 4224 0 11 23 0 0 4
404 213
518 213
518 242
602 242
1 6 18 0 0 4224 0 13 23 0 0 4
404 187
537 187
537 233
602 233
1 5 19 0 0 4224 0 14 23 0 0 4
404 161
556 161
556 224
602 224
19 1 20 0 0 8320 0 23 22 0 0 3
678 260
700 260
700 301
20 1 21 0 0 4224 0 23 21 0 0 3
678 269
733 269
733 301
21 1 22 0 0 4224 0 23 20 0 0 3
678 278
765 278
765 301
22 1 23 0 0 4224 0 23 19 0 0 3
678 287
798 287
798 301
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
